module MD5Controller(
    input clock,
    input [2:0] increment,
    input [7:0] startingPosition,
    input [127:0] target_hash,
    output reg hashes_equal,
    output [127:0] reg plaintext
);



endmodule